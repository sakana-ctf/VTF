module vlog

import term

pub const false_log = term.red('[False] ')
pub const true_log = term.green('[True] ')
pub const set_log = term.yellow('[Setting] ')
pub const warn_log = term.yellow('[Warn] ')
pub const threat_log = term.red('[Threat] ')




